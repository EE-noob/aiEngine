`ifndef ics_mem_model_PKG_SV
`define ics_mem_model_PKG_SV


package ics_mem_model_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    `include "ics_mem_model.sv"

endpackage: ics_mem_model_pkg

`endif

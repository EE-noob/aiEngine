`ifndef ics_monitor_PKG_SV
`define ics_monitor_PKG_SV


package ics_monitor_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    `include "ics_monitor.sv"

endpackage: ics_monitor_pkg

`endif

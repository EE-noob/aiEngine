// case209_define.vh  –  Auto-gen by ics_testgen.py

`define ICS_INPUT_DATA       "../../data/ics_input_data7.txt"
`define ICS_INTLV_OUT_DATA   "../../data/ics_intlv_out_data7.txt"
`define ICS_OUTPUT_DATA      "../../data/ics_output_data7.txt"
`define ICS_SCRAMBLE_CODE    "../../data/ics_scram_code7.txt"

`define GROUP_WIDTH_ARRAY_0 \
  '{ 6, 6, 5, 5, 4, 3, 2, 1 }
`define GROUP_WIDTH_ARRAY_1 \
  '{ 6, 6, 5, 5, 4, 3, 2, 1 }
`define GROUP_WIDTH_ARRAY_2 \
  '{ 6, 6, 5, 5, 4, 3, 2, 1 }
`define GOLDEN_LINES_PER_PART '{1, 1, 1}
`define ICS_SCRAMBLE_OUTPUT_NUM 1

`define ICS_C_INIT             31'h11
`define ICS_Q_SIZE             4'd2
`define ICS_PART0_EN           1'b1
`define ICS_PART0_N_SIZE       11'd32
`define ICS_PART0_E_SIZE       14'd32
`define ICS_PART0_L_SIZE       14'd2
`define ICS_PART0_ST_IDX       14'd31
`define ICS_PART1_EN           1'b1
`define ICS_PART1_N_SIZE       11'd32
`define ICS_PART1_E_SIZE       14'd32
`define ICS_PART1_L_SIZE       14'd2
`define ICS_PART1_ST_IDX       14'd31
`define ICS_PART2_EN           1'b1
`define ICS_PART2_N_SIZE       11'd32
`define ICS_PART2_E_SIZE       14'd32
`define ICS_PART2_L_SIZE       14'd2
`define ICS_PART2_ST_IDX       14'd31

`ifndef ics_mst_PKG_SV
`define ics_mst_PKG_SV


package ics_mst_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    
    `include "ics_mst_agent_cfg_base.sv"
    `include "ics_mst_agent_cfg.sv"
    `include "ics_mst_tr.sv"
    `include "ics_mst_coverage.sv"
    `include "ics_mst_sequencer.sv"
    `include "ics_mst_monitor.sv"
    `include "ics_mst_driver.sv"
    `include "ics_mst_reg_adapter.sv"
    `include "ics_mst_agent.sv"

endpackage: ics_mst_pkg

`endif

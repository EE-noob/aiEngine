`ifndef combine_checker_PKG_SV
`define combine_checker_PKG_SV


package combine_checker_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    `include "combine_checker.sv"

endpackage: combine_checker_pkg

`endif

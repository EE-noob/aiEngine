`ifndef filo_collector_PKG_SV
`define filo_collector_PKG_SV


package filo_collector_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;
    `include "filo_collector.sv"

endpackage: filo_collector_pkg

`endif
